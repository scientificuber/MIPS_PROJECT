module main()

endmodule;
