module instruction_memory(address,data_out);
input [31:0]address;
output  [31:0] data_out;
reg [31:0]memory[360:0];
initial begin

		//load word t0 512(s0)
		memory[0]=32'b100011_01000_10000_0000001000000000;
		//load word t1 768(s0)
		memory[4]=32'b100011_01001_10000_0000001100000000;
		//load word t2 516(s0)
		memory[8]=32'b100011_01010_10000_0000001000000100;
		//load word t3 772(s0)
		memory[12]=32'b100011_01011_10000_0000001100000100;
		//load word t4 520(s0)
		memory[16]=32'b100011_01100_10000_0000001000001000;
		//load word t5 776(s0)
		memory[20]=32'b100011_01101_10000_0000001100001000;
		//mul t6 t0 t1
		memory[24]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[28]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[32]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[36]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[40]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store word t6 256(s0)
		memory[44]=33'b101011_01110_10000_0000000100000000;
		//
		// /*
		//load word t1 780(s0)
		memory[48]=32'b100011_01001_10000_0000001100001100;
		//load word t3 784(s0)
		memory[52]=32'b100011_01011_10000_0000001100010000;
		//load word t5 788(s0)
		memory[56]=32'b100011_01101_10000_0000001100010100;
		//mul t6 t0 t1
		memory[60]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[64]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[68]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[72]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[76]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store word t6 260(s0)
		memory[80]=32'b101011_01110_10000_0000000100000100;
		//
		//load word t1 792(s0)
		memory[84]=32'b100011_01001_10000_0000001100011000;
		//load word t3 796(s0)
		memory[88]=32'b100011_01011_10000_0000001100011100;
		//load word t5 800(s0)
		memory[92]=32'b100011_01101_10000_0000001100100000;
		//mul t6 t0 t1
		memory[96]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[100]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[104]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[108]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[112]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store word t6 264(s0)
		memory[116]=32'b101011_01110_10000_0000000100001000;
		//
		//load word t0 524(s0)
		memory[120]=32'b100011_01000_10000_0000001000001100;
		//load word t2 528(s0)
		memory[124]=32'b100011_01010_10000_0000001000010000;
		//load word t4 532(s0)
		memory[128]=32'b100011_01100_10000_0000001000010100;
		//load word t1 768(s0)
		memory[132]=32'b100011_01001_10000_0000001100000000;
		//load word t3 772(s0)
		memory[136]=32'b100011_01011_10000_0000001100000100;
		//load word t5 776(s0)
		memory[140]=32'b100011_01101_10000_0000001100001000;
		//mul t6 t0 t1
		memory[144]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[148]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[152]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[156]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[160]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store word t6 268(s0)
		memory[164]=32'b101011_01110_10000_0000000100001100;
		//
		//load t1 780(s0)
		memory[168]=32'b100011_01001_10000_0000001100001100;
		//load t3 784(s0)
		memory[172]=32'b100011_01011_10000_0000001100010000;
		//load t5 788(s0)
		memory[176]=32'b100011_01101_10000_0000001100010100;
		//mul t6 t0 t1
		memory[180]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[184]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[188]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[192]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[196]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store word t6 272(s0)
		memory[200]=32'b101011_01110_10000_0000000100010000;
		//
		//load t1 792(s0)
		memory[204]=32'b100011_01001_10000_0000001100011000;
		//load t3 796(s0)
		memory[208]=32'b100011_01011_10000_0000001100011100;
		//load t5 800(s0)
		memory[212]=32'b100011_01101_10000_0000001100100000;
		//mul t6 t0 t1
		memory[216]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[220]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[224]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[228]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[232]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store word t6 276(s0)
		memory[236]=32'b101011_01110_10000_0000000100010100;
		//
		//load t0 536(s0)
		memory[240]=32'b100011_01000_10000_0000001000011000;
		//load t2 540(s0)
		memory[244]=32'b100011_01010_10000_0000001000011100;
		//load t4 544(s0)
		memory[248]=32'b100011_01100_10000_0000001000100000;
		//load t1 768(s0)
		memory[252]=32'b100011_01001_10000_0000001100000000;
		//load t3 772(s0)
		memory[256]=32'b100011_01011_10000_0000001100000100;
		//load t5 776(s0)
		memory[260]=32'b100011_01101_10000_0000001100001000;
		//mul t6 t0 t1
		memory[264]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[268]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[272]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[276]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[280]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store word t6 280(s0)
		memory[284]=32'b101011_01110_10000_0000000100011000;
		//
		//load t1 780(s0)
		memory[288]=32'b100011_01001_10000_0000001100001100;
		//load t3 784(s0)
		memory[292]=32'b100011_01011_10000_0000001100010000;
		//load t5 788(s0)
		memory[296]=32'b100011_01101_10000_0000001100010100;
		//mul t6 t0 t1
		memory[300]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[304]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[308]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[312]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[316]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store t6 284(s0)
		memory[320]=32'b101011_01110_10000_0000000100011100;
		//
		//load t1 792(s0)
		memory[324]=32'b100011_01001_10000_0000001100011000;
		//load t3 796(s0)
		memory[328]=32'b100011_01011_10000_0000001100011100;
		//load t5 800(s0)
		memory[332]=32'b100011_01101_10000_0000001100100000;
		//mul t6 t0 t1
		memory[336]=32'b000000_01110_01000_01001_00000_011000;
		//mul t7 t2 t3
		memory[340]=32'b000000_01111_01010_01011_00000_011000;
		//mul s5 t4 t5
		memory[344]=32'b000000_10101_01100_01101_00000_011000;
		//add t6 t6 t7
		memory[348]=32'b000000_01110_01110_01111_00000_100000;
		//add t6 t6 s5
		memory[352]=32'b000000_01110_01110_10101_00000_100000;
		//
		//store t6 288(s0)
		memory[356]=32'b101011_01110_10000_0000000100100000;
		//
		// */
end
assign data_out=memory[address];
// always @ ( * ) begin
// 	data_out = memory[address];
// 	$display("%b", data_out);
// end
endmodule
